// %u %z
